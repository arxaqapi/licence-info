LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TP1EX1 IS
	PORT (  E2, E1, E0		: IN STD_LOGIC;
		S3, S2, S1, S0	: OUT STD_LOGIC);
END ENTITY TP1EX1;

ARCHITECTURE fdd_TP1EX1 OF TP1EX1 IS
	SIGNAL S : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SUBTYPE selecteur IS STD_LOGIC_VECTOR(2 DOWNTO 0);
BEGIN
	(S3, S2, S1, S0) <= S;
	WITH selecteur'( E2 & E1 & E0 ) SELECT
		S <=	"0001" WHEN "000",
			"0010" WHEN "001",
			"0100" WHEN "010",
			"1000" WHEN "011",
			"ZZZZ" WHEN "100",
			"ZZZZ" WHEN "101",
			"ZZZZ" WHEN "110",
			"ZZZZ" WHEN "111",
			"0000" WHEN OTHERS;
END ARCHITECTURE fdd_TP1EX1;
