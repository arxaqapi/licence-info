LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ADD1B IS
	PORT (  a, b, c	: IN STD_LOGIC;
		S, R	: OUT STD_LOGIC);
END ENTITY ADD1B;

ARCHITECTURE fdd_ADD1B OF ADD1B IS
	SIGNAL SORT : STD_LOGIC_VECTOR(1 DOWNTO 0);
	SUBTYPE selecteur IS STD_LOGIC_VECTOR(2 DOWNTO 0);
BEGIN
	(S, R) <= SORT;
	WITH selecteur'( a & b & c ) SELECT
		SORT <=	"00" WHEN "000",
			"10" WHEN "001",
			"10" WHEN "010",
			"01" WHEN "011",
			"10" WHEN "100",
			"01" WHEN "101",
			"01" WHEN "110",
			"11" WHEN "111",
			"00" WHEN OTHERS;
END ARCHITECTURE fdd_ADD1B;
